module hello_tb;

    initial begin
        $display("Hello, System Verilog!");
        $stop;
    end
    
endmodule