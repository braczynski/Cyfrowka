module not1 (
        output logic y,
        input logic a
);

assign y = ~a;

endmodule

