module nor2 (
        output logic y,
        input logic a,
        input logic b
);

assign y = ~(a | b);

endmodule

